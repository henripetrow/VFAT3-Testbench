------------------------------------------------------------------------------
--   ____  ____
--  /   /\/   /
-- /___/  \  /    Vendor: Xilinx
-- \   \   \/     Version : 2.1
--  \   \         Application : 7 Series FPGAs Transceivers Wizard 
--  /   /         Filename : gig_eth_pcs_pma_v11_4_gtwizard_init.vhd
-- /___/   /\      
-- \   \  /  \ 
--  \___\/\___\
--
--  Description : This module instantiates the modules required for
--                reset and initialisation of the Transceiver
--
-- Module GTWIZARD_init
-- Generated by Xilinx 7 Series FPGAs Transceivers Wizard
-- 
-- 
-- (c) Copyright 2010-2012 Xilinx, Inc. All rights reserved.
-- 
-- This file contains confidential and proprietary information
-- of Xilinx, Inc. and is protected under U.S. and
-- international copyright and other intellectual property
-- laws.
-- 
-- DISCLAIMER
-- This disclaimer is not a license and does not grant any
-- rights to the materials distributed herewith. Except as
-- otherwise provided in a valid license issued to you by
-- Xilinx, and to the maximum extent permitted by applicable
-- law: (1) THESE MATERIALS ARE MADE AVAILABLE "AS IS" AND
-- WITH ALL FAULTS, AND XILINX HEREBY DISCLAIMS ALL WARRANTIES
-- AND CONDITIONS, EXPRESS, IMPLIED, OR STATUTORY, INCLUDING
-- BUT NOT LIMITED TO WARRANTIES OF MERCHANTABILITY, NON-
-- INFRINGEMENT, OR FITNESS FOR ANY PARTICULAR PURPOSE; and
-- (2) Xilinx shall not be liable (whether in contract or tort,
-- including negligence, or under any other theory of
-- liability) for any loss or damage of any kind or nature
-- related to, arising under or in connection with these
-- materials, including for any direct, or any indirect,
-- special, incidental, or consequential loss or damage
-- (including loss of data, profits, goodwill, or any type of
-- loss or damage suffered as a result of any action brought
-- by a third party) even if such damage or loss was
-- reasonably foreseeable or Xilinx had been advised of the
-- possibility of the same.
-- 
-- CRITICAL APPLICATIONS
-- Xilinx products are not designed or intended to be fail-
-- safe, or for use in any application requiring fail-safe
-- performance, such as life-support or safety devices or
-- systems, Class III medical devices, nuclear facilities,
-- applications related to the deployment of airbags, or any
-- other applications that could lead to death, personal
-- injury, or severe property or environmental damage
-- (individually and collectively, "Critical
-- Applications"). Customer assumes the sole risk and
-- liability of any use of Xilinx products in Critical
-- Applications, subject only to applicable laws and
-- regulations governing limitations on product liability.
-- 
-- THIS COPYRIGHT NOTICE AND DISCLAIMER MUST BE RETAINED AS
-- PART OF THIS FILE AT ALL TIMES. 


library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use ieee.std_logic_unsigned.all;
library UNISIM;
use UNISIM.VCOMPONENTS.ALL;

--***********************************Entity Declaration************************

entity gig_eth_pcs_pma_v11_4_GTWIZARD_init is
generic
(
    EXAMPLE_SIM_GTRESET_SPEEDUP             : string    := "TRUE";     -- simulation setting for GT SecureIP model
    EXAMPLE_SIMULATION                      : integer   := 0;          -- Set to 1 for simulation
    EXAMPLE_USE_CHIPSCOPE                   : integer   := 0           -- Set to 1 to use Chipscope to drive resets

);
port
(
    SYSCLK_IN                               : in   std_logic;
    SOFT_RESET_IN                           : in   std_logic;
    GT0_TX_FSM_RESET_DONE_OUT               : out  std_logic;
    GT0_RX_FSM_RESET_DONE_OUT               : out  std_logic;
    GT0_DATA_VALID_IN                       : in   std_logic;

    --_________________________________________________________________________
    --GT0  (X1Y4)
    --____________________________CHANNEL PORTS________________________________
    ------------------------- Channel - Ref Clock Ports ------------------------
    GT0_GTREFCLK0_IN                        : in   std_logic;
    -------------------------------- Channel PLL -------------------------------
    GT0_CPLLFBCLKLOST_OUT                   : out  std_logic;
    GT0_CPLLLOCK_OUT                        : out  std_logic;
    GT0_CPLLLOCKDETCLK_IN                   : in   std_logic;
    GT0_CPLLRESET_IN                        : in   std_logic;
    ------------------------------- Eye Scan Ports -----------------------------
    GT0_EYESCANDATAERROR_OUT                : out  std_logic;
    ------------------------ Loopback and Powerdown Ports ----------------------
    GT0_LOOPBACK_IN                         : in   std_logic_vector(2 downto 0);
    GT0_RXPD_IN                             : in   std_logic_vector(1 downto 0);
    GT0_TXPD_IN                             : in   std_logic_vector(1 downto 0);
    ------------------------------- Receive Ports ------------------------------
    GT0_RXUSERRDY_IN                        : in   std_logic;
    ----------------------- Receive Ports - 8b10b Decoder ----------------------
    GT0_RXCHARISCOMMA_OUT                   : out  std_logic_vector(1 downto 0);
    GT0_RXCHARISK_OUT                       : out  std_logic_vector(1 downto 0);
    GT0_RXDISPERR_OUT                       : out  std_logic_vector(1 downto 0);
    GT0_RXNOTINTABLE_OUT                    : out  std_logic_vector(1 downto 0);
    ------------------- Receive Ports - Clock Correction Ports -----------------
        GT0_RXCLKCORCNT_OUT                     : out  std_logic_vector(1 downto 0);
        --------------- Receive Ports - Comma Detection and Alignment --------------
    GT0_RXMCOMMAALIGNEN_IN                  : in   std_logic;
    GT0_RXPCOMMAALIGNEN_IN                  : in   std_logic;
    ------------------- Receive Ports - RX Data Path interface -----------------
    GT0_GTRXRESET_IN                        : in   std_logic;
    GT0_RXDATA_OUT                          : out  std_logic_vector(15 downto 0);
    GT0_RXOUTCLK_OUT                        : out  std_logic;
    GT0_RXUSRCLK_IN                         : in   std_logic;
    GT0_RXUSRCLK2_IN                        : in   std_logic;
    ------- Receive Ports - RX Driver,OOB signalling,Coupling and Eq.,CDR ------
    GT0_GTXRXN_IN                           : in   std_logic;
    GT0_GTXRXP_IN                           : in   std_logic;
    GT0_RXCDRLOCK_OUT                       : out  std_logic;
    GT0_RXELECIDLE_OUT                      : out  std_logic;
    -------- Receive Ports - RX Elastic Buffer and Phase Alignment Ports -------
    GT0_RXBUFRESET_IN                       : in   std_logic;
    GT0_RXBUFSTATUS_OUT                     : out  std_logic_vector(2 downto 0);
    ------------------------ Receive Ports - RX PLL Ports ----------------------
    GT0_RXRESETDONE_OUT                     : out  std_logic;
    ------------------------------- Transmit Ports -----------------------------
    GT0_TXUSERRDY_IN                        : in   std_logic;
    ---------------- Transmit Ports - 8b10b Encoder Control Ports --------------
    GT0_TXCHARDISPMODE_IN                   : in   std_logic_vector(1 downto 0);
    GT0_TXCHARDISPVAL_IN                    : in   std_logic_vector(1 downto 0);
    GT0_TXCHARISK_IN                        : in   std_logic_vector(1 downto 0);
    ------------ Transmit Ports - TX Buffer and Phase Alignment Ports ----------
    GT0_TXBUFSTATUS_OUT                     : out  std_logic_vector(1 downto 0);
    ------------------ Transmit Ports - TX Data Path interface -----------------
    GT0_GTTXRESET_IN                        : in   std_logic;
    GT0_TXDATA_IN                           : in   std_logic_vector(15 downto 0);
    GT0_TXOUTCLK_OUT                        : out  std_logic;
    GT0_TXOUTCLKFABRIC_OUT                  : out  std_logic;
    GT0_TXOUTCLKPCS_OUT                     : out  std_logic;
    GT0_TXUSRCLK_IN                         : in   std_logic;
    GT0_TXUSRCLK2_IN                        : in   std_logic;
    ---------------- Transmit Ports - TX Driver and OOB signaling --------------
    GT0_GTXTXN_OUT                          : out  std_logic;
    GT0_GTXTXP_OUT                          : out  std_logic;
    ----------------------- Transmit Ports - TX PLL Ports ----------------------
    GT0_TXRESETDONE_OUT                     : out  std_logic



);

end gig_eth_pcs_pma_v11_4_GTWIZARD_init;
    
architecture RTL of gig_eth_pcs_pma_v11_4_GTWIZARD_init is

--**************************Component Declarations*****************************


component gig_eth_pcs_pma_v11_4_GTWIZARD 
generic
(
    -- Simulation attributes
    WRAPPER_SIM_GTRESET_SPEEDUP    : string    := "FALSE" -- Set to 1 to speed up sim reset

);
port
(

    --_________________________________________________________________________
    --_________________________________________________________________________
    --GT0  (X1Y4)
    --____________________________CHANNEL PORTS________________________________
    ------------------------- Channel - Ref Clock Ports ------------------------
    GT0_GTREFCLK0_IN                        : in   std_logic;
    -------------------------------- Channel PLL -------------------------------
    GT0_CPLLFBCLKLOST_OUT                   : out  std_logic;
    GT0_CPLLLOCK_OUT                        : out  std_logic;
    GT0_CPLLLOCKDETCLK_IN                   : in   std_logic;
    GT0_CPLLREFCLKLOST_OUT                  : out  std_logic;
    GT0_CPLLRESET_IN                        : in   std_logic;
    ------------------------------- Eye Scan Ports -----------------------------
    GT0_EYESCANDATAERROR_OUT                : out  std_logic;
    ------------------------ Loopback and Powerdown Ports ----------------------
    GT0_LOOPBACK_IN                         : in   std_logic_vector(2 downto 0);
    GT0_RXPD_IN                             : in   std_logic_vector(1 downto 0);
    GT0_TXPD_IN                             : in   std_logic_vector(1 downto 0);
    ------------------------------- Receive Ports ------------------------------
    GT0_RXUSERRDY_IN                        : in   std_logic;
    ----------------------- Receive Ports - 8b10b Decoder ----------------------
    GT0_RXCHARISCOMMA_OUT                   : out  std_logic_vector(1 downto 0);
    GT0_RXCHARISK_OUT                       : out  std_logic_vector(1 downto 0);
    GT0_RXDISPERR_OUT                       : out  std_logic_vector(1 downto 0);
    GT0_RXNOTINTABLE_OUT                    : out  std_logic_vector(1 downto 0);
    ------------------- Receive Ports - Clock Correction Ports -----------------
        GT0_RXCLKCORCNT_OUT                     : out  std_logic_vector(1 downto 0);
        --------------- Receive Ports - Comma Detection and Alignment --------------
    GT0_RXMCOMMAALIGNEN_IN                  : in   std_logic;
    GT0_RXPCOMMAALIGNEN_IN                  : in   std_logic;
    ------------------- Receive Ports - RX Data Path interface -----------------
    GT0_GTRXRESET_IN                        : in   std_logic;
    GT0_RXDATA_OUT                          : out  std_logic_vector(15 downto 0);
    GT0_RXOUTCLK_OUT                        : out  std_logic;
    GT0_RXPCSRESET_IN                       : in   std_logic;
    GT0_RXUSRCLK_IN                         : in   std_logic;
    GT0_RXUSRCLK2_IN                        : in   std_logic;
    ------- Receive Ports - RX Driver,OOB signalling,Coupling and Eq.,CDR ------
    GT0_GTXRXN_IN                           : in   std_logic;
    GT0_GTXRXP_IN                           : in   std_logic;
    GT0_RXCDRLOCK_OUT                       : out  std_logic;
    GT0_RXELECIDLE_OUT                      : out  std_logic;
    -------- Receive Ports - RX Elastic Buffer and Phase Alignment Ports -------
    GT0_RXBUFRESET_IN                       : in   std_logic;
    GT0_RXBUFSTATUS_OUT                     : out  std_logic_vector(2 downto 0);
    ------------------------ Receive Ports - RX PLL Ports ----------------------
    GT0_RXRESETDONE_OUT                     : out  std_logic;
    ------------------------------- Transmit Ports -----------------------------
    GT0_TXUSERRDY_IN                        : in   std_logic;
    ---------------- Transmit Ports - 8b10b Encoder Control Ports --------------
    GT0_TXCHARDISPMODE_IN                   : in   std_logic_vector(1 downto 0);
    GT0_TXCHARDISPVAL_IN                    : in   std_logic_vector(1 downto 0);
    GT0_TXCHARISK_IN                        : in   std_logic_vector(1 downto 0);
    ------------ Transmit Ports - TX Buffer and Phase Alignment Ports ----------
    GT0_TXBUFSTATUS_OUT                     : out  std_logic_vector(1 downto 0);
    ------------------ Transmit Ports - TX Data Path interface -----------------
    GT0_GTTXRESET_IN                        : in   std_logic;
    GT0_TXDATA_IN                           : in   std_logic_vector(15 downto 0);
    GT0_TXOUTCLK_OUT                        : out  std_logic;
    GT0_TXOUTCLKFABRIC_OUT                  : out  std_logic;
    GT0_TXOUTCLKPCS_OUT                     : out  std_logic;
    GT0_TXPCSRESET_IN                       : in   std_logic;
    GT0_TXUSRCLK_IN                         : in   std_logic;
    GT0_TXUSRCLK2_IN                        : in   std_logic;
    ---------------- Transmit Ports - TX Driver and OOB signaling --------------
    GT0_GTXTXN_OUT                          : out  std_logic;
    GT0_GTXTXP_OUT                          : out  std_logic;
    ----------------------- Transmit Ports - TX PLL Ports ----------------------
    GT0_TXRESETDONE_OUT                     : out  std_logic
   


);
end component;

component gig_eth_pcs_pma_v11_4_TX_STARTUP_FSM
  Generic(
           GT_TYPE                  : string := "GTX";
           STABLE_CLOCK_PERIOD      : integer range 4 to 20 := 8; --Period of the stable clock driving this state-machine, unit is [ns]
           RETRY_COUNTER_BITWIDTH   : integer range 2 to 8  := 8; 
            TX_QPLL_USED             : boolean := False;           -- the TX and RX Reset FSMs must
           RX_QPLL_USED             : boolean := False;           -- share these two generic values
           PHASE_ALIGNMENT_MANUAL   : boolean := True             -- Decision if a manual phase-alignment is necessary or the automatic 
                                                                  -- is enough. For single-lane applications the automatic alignment is 
                                                                  -- sufficient              
         );     
    Port ( STABLE_CLOCK             : in  STD_LOGIC;              --Stable Clock, either a stable clock from the PCB
                                                                  --or reference-clock present at startup.
           TXUSERCLK                : in  STD_LOGIC;              --TXUSERCLK as used in the design
           SOFT_RESET               : in  STD_LOGIC;              --User Reset, can be pulled any time
           QPLLREFCLKLOST           : in  STD_LOGIC;              --QPLL Reference-clock for the GT is lost
           CPLLREFCLKLOST           : in  STD_LOGIC;              --CPLL Reference-clock for the GT is lost
           QPLLLOCK                 : in  STD_LOGIC;              --Lock Detect from the QPLL of the GT
           CPLLLOCK                 : in  STD_LOGIC;              --Lock Detect from the CPLL of the GT
           TXRESETDONE              : in  STD_LOGIC;      
           MMCM_LOCK                : in  STD_LOGIC;      
           GTTXRESET                : out STD_LOGIC:='0';      
           MMCM_RESET               : out STD_LOGIC:='0';      
           QPLL_RESET               : out STD_LOGIC:='0';        --Reset QPLL
           CPLL_RESET               : out STD_LOGIC:='0';        --Reset CPLL
           TX_FSM_RESET_DONE        : out STD_LOGIC:='0';        --Reset-sequence has sucessfully been finished.
           TXUSERRDY                : out STD_LOGIC:='0';
           RUN_PHALIGNMENT          : out STD_LOGIC:='0';
           RESET_PHALIGNMENT        : out STD_LOGIC:='0';
           PHALIGNMENT_DONE         : in  STD_LOGIC;
           
           RETRY_COUNTER            : out  STD_LOGIC_VECTOR (RETRY_COUNTER_BITWIDTH-1 downto 0):=(others=>'0')-- Number of 
                                                            -- Retries it took to get the transceiver up and running
           );
end component;

component gig_eth_pcs_pma_v11_4_RX_STARTUP_FSM
  Generic(
           EXAMPLE_SIMULATION       : integer := 0;
           EQ_MODE                  : string := "DFE";
           GT_TYPE                  : string := "GTX";
           STABLE_CLOCK_PERIOD      : integer range 4 to 20 := 8; --Period of the stable clock driving this state-machine, unit is [ns]
           RETRY_COUNTER_BITWIDTH   : integer range 2 to 8  := 8; 
           TX_QPLL_USED             : boolean := False;           -- the TX and RX Reset FSMs must
           RX_QPLL_USED             : boolean := False;           -- share these two generic values
           PHASE_ALIGNMENT_MANUAL   : boolean := True             -- Decision if a manual phase-alignment is necessary or the automatic 
                                                                  -- is enough. For single-lane applications the automatic alignment is 
                                                                  -- sufficient                         
         );     
    Port ( STABLE_CLOCK             : in  STD_LOGIC;        --Stable Clock, either a stable clock from the PCB
                                                            --or reference-clock present at startup.
           RXUSERCLK                : in  STD_LOGIC;        --RXUSERCLK as used in the design
           SOFT_RESET               : in  STD_LOGIC;        --User Reset, can be pulled any time
           QPLLREFCLKLOST           : in  STD_LOGIC;        --QPLL Reference-clock for the GT is lost
           CPLLREFCLKLOST           : in  STD_LOGIC;        --CPLL Reference-clock for the GT is lost
           QPLLLOCK                 : in  STD_LOGIC;        --Lock Detect from the QPLL of the GT
           CPLLLOCK                 : in  STD_LOGIC;        --Lock Detect from the CPLL of the GT
           RXRESETDONE              : in  STD_LOGIC;
           MMCM_LOCK                : in  STD_LOGIC;
           RECCLK_STABLE            : in  STD_LOGIC;
           RECCLK_MONITOR_RESTART   : in  STD_LOGIC;
           DATA_VALID               : in  STD_LOGIC;
           TXUSERRDY                : in  STD_LOGIC;       --TXUSERRDY from GT 
           GTRXRESET                : out STD_LOGIC:='0';
           MMCM_RESET               : out STD_LOGIC:='0';
           QPLL_RESET               : out STD_LOGIC:='0';  --Reset QPLL (only if RX uses QPLL)
           CPLL_RESET               : out STD_LOGIC:='0';  --Reset CPLL (only if RX uses CPLL)
           RX_FSM_RESET_DONE        : out STD_LOGIC:='0';  --Reset-sequence has sucessfully been finished.
           RXUSERRDY                : out STD_LOGIC:='0';
           RUN_PHALIGNMENT          : out STD_LOGIC;
           PHALIGNMENT_DONE         : in  STD_LOGIC; 
           RESET_PHALIGNMENT        : out STD_LOGIC:='0';           
           RXDFEAGCHOLD             : out STD_LOGIC;
           RXDFELFHOLD              : out STD_LOGIC;
           RXLPMLFHOLD              : out STD_LOGIC;
           RXLPMHFHOLD              : out STD_LOGIC;
           RETRY_COUNTER            : out STD_LOGIC_VECTOR (RETRY_COUNTER_BITWIDTH-1 downto 0):=(others=>'0')-- Number of 
                                                            -- Retries it took to get the transceiver up and running
           );
end component;

--**************************Component Declarations*****************************

component gig_eth_pcs_pma_v11_4_sync_block
generic (
  INITIALISE : bit_vector(1 downto 0) := "00"
);
port  (
          clk           : in  std_logic;
          data_in       : in  std_logic;
          data_out      : out std_logic
       );
end component;

  function get_cdrlock_time(is_sim : in integer) return integer is
    variable lock_time: integer;
  begin
    if (is_sim = 1) then
      lock_time := 1000;
    else
      lock_time := 50000 / integer(1.25); --Typical CDR lock time is 50,000UI as per DS183
    end if;
    return lock_time;
  end function;

--***********************************Parameter Declarations********************

    constant DLY : time := 1 ns;
    constant STABLE_CLOCK_PERIOD  : integer := 5;  --Period of the stable clock driving this state-machine, unit is [ns]
    constant RX_CDRLOCK_TIME      : integer := get_cdrlock_time(EXAMPLE_SIMULATION);       -- 200us
    constant WAIT_TIME_CDRLOCK    : integer := RX_CDRLOCK_TIME / STABLE_CLOCK_PERIOD;      -- 200 us time-out

    -------------------------- GT Wrapper Wires ------------------------------
    signal   gt0_cpllreset_i                 : std_logic;
    signal   gt0_cpllreset_t                 : std_logic;
    signal   gt0_cpllrefclklost_i            : std_logic;
    signal   gt0_cplllock_i                  : std_logic;
    signal   gt0_txresetdone_i               : std_logic;
    signal   gt0_rxresetdone_i               : std_logic;
    signal   gt0_gttxreset_i                 : std_logic;
    signal   gt0_gttxreset_t                 : std_logic;
    signal   gt0_gtrxreset_i                 : std_logic;
    signal   gt0_gtrxreset_t                 : std_logic;
    signal   gt0_txpcsreset_i                : std_logic;
    signal   gt0_rxpcsreset_i                : std_logic;
    signal   gt0_txuserrdy_i                 : std_logic;
    signal   gt0_txuserrdy_t                 : std_logic;
    signal   gt0_rxuserrdy_i                 : std_logic;
    signal   gt0_rxuserrdy_t                 : std_logic;

    signal   gt0_rxdfeagchold_i              : std_logic;
    signal   gt0_rxdfelfhold_i               : std_logic;
    signal   gt0_rxlpmlfhold_i               : std_logic;
    signal   gt0_rxlpmhfhold_i               : std_logic;

    ------------------------------- Global Signals -----------------------------
    signal  tied_to_ground_i                : std_logic;
    signal  tied_to_vcc_i                   : std_logic;

    signal   gt0_rxoutclk_i                  : std_logic;
    signal   gt0_recclk_stable_i             : std_logic;
    signal   gt0_rxelecidle_i                : std_logic;

    signal   rx_cdrlock_counter  :   integer range 0 to WAIT_TIME_CDRLOCK:= 0 ;
    signal      rx_cdrlocked                    : std_logic;

    signal   gt0_txresetdone_sync            : std_logic;
    signal   gt0_rxresetdone_sync            : std_logic;
    signal   gt0_gtrxreset_gt                : std_logic;
    signal   gt0_gttxreset_gt                : std_logic;
--**************************** Main Body of Code *******************************
begin
    --  Static signal Assigments
    tied_to_ground_i                             <= '0';
    tied_to_vcc_i                                <= '1';
    gt0_cpllrefclklost_i <= '0';
   gt0_gttxreset_gt                             <= gt0_gttxreset_t or GT0_GTTXRESET_IN; 
    gt0_gtrxreset_gt                             <= gt0_gtrxreset_t or GT0_GTRXRESET_IN; 

sync_block_txresetdone : gig_eth_pcs_pma_v11_4_sync_block 
  port map (
             clk             => SYSCLK_IN,
             data_in         => gt0_txresetdone_i,
             data_out        => gt0_txresetdone_sync
          );

sync_block_rxresetdone : gig_eth_pcs_pma_v11_4_sync_block 
  port map (
             clk             => SYSCLK_IN,
             data_in         => gt0_rxresetdone_i,
             data_out        => gt0_rxresetdone_sync
          );
    ----------------------------- The GT Wrapper -----------------------------
    
    -- Use the instantiation template in the example directory to add the GT wrapper to your design.
    -- In this example, the wrapper is wired up for basic operation with a frame generator and frame 
    -- checker. The GTs will reset, then attempt to align and transmit data. If channel bonding is 
    -- enabled, bonding should occur after alignment.


    GTWIZARD_i : gig_eth_pcs_pma_v11_4_GTWIZARD
    generic map
    (
        WRAPPER_SIM_GTRESET_SPEEDUP     =>      EXAMPLE_SIM_GTRESET_SPEEDUP
    )
    port map
    (
  
        --_____________________________________________________________________
        --_____________________________________________________________________
        --GT0  (X1Y4)

        ------------------------- Channel - Ref Clock Ports ------------------------
        GT0_GTREFCLK0_IN                =>      GT0_GTREFCLK0_IN,
        -------------------------------- Channel PLL -------------------------------
        GT0_CPLLFBCLKLOST_OUT           =>      GT0_CPLLFBCLKLOST_OUT,
        GT0_CPLLLOCK_OUT                =>      gt0_cplllock_i,
        GT0_CPLLLOCKDETCLK_IN           =>      GT0_CPLLLOCKDETCLK_IN,
        GT0_CPLLREFCLKLOST_OUT          =>      open,
        GT0_CPLLRESET_IN                =>      gt0_cpllreset_i,
        ------------------------------- Eye Scan Ports -----------------------------
        GT0_EYESCANDATAERROR_OUT        =>      GT0_EYESCANDATAERROR_OUT,
        ------------------------ Loopback and Powerdown Ports ----------------------
        GT0_LOOPBACK_IN                 =>      GT0_LOOPBACK_IN,
        GT0_RXPD_IN                     =>      GT0_RXPD_IN,
        GT0_TXPD_IN                     =>      GT0_TXPD_IN,
        ------------------------------- Receive Ports ------------------------------
        GT0_RXUSERRDY_IN                =>      gt0_rxuserrdy_i,
        ----------------------- Receive Ports - 8b10b Decoder ----------------------
        GT0_RXCHARISCOMMA_OUT           =>      GT0_RXCHARISCOMMA_OUT,
        GT0_RXCHARISK_OUT               =>      GT0_RXCHARISK_OUT,
        GT0_RXDISPERR_OUT               =>      GT0_RXDISPERR_OUT,
        GT0_RXNOTINTABLE_OUT            =>      GT0_RXNOTINTABLE_OUT,
        ------------------- Receive Ports - Clock Correction Ports -----------------
                GT0_RXCLKCORCNT_OUT             =>      GT0_RXCLKCORCNT_OUT,
                --------------- Receive Ports - Comma Detection and Alignment --------------
        GT0_RXMCOMMAALIGNEN_IN          =>      GT0_RXMCOMMAALIGNEN_IN,
        GT0_RXPCOMMAALIGNEN_IN          =>      GT0_RXPCOMMAALIGNEN_IN,
        ------------------- Receive Ports - RX Data Path interface -----------------
        GT0_GTRXRESET_IN                =>      gt0_gtrxreset_gt,
        GT0_RXDATA_OUT                  =>      GT0_RXDATA_OUT,
        GT0_RXOUTCLK_OUT                =>      gt0_rxoutclk_i,
        GT0_RXPCSRESET_IN               =>      gt0_rxpcsreset_i,
        GT0_RXUSRCLK_IN                 =>      GT0_RXUSRCLK_IN,
        GT0_RXUSRCLK2_IN                =>      GT0_RXUSRCLK2_IN,
        ------- Receive Ports - RX Driver,OOB signalling,Coupling and Eq.,CDR ------
        GT0_GTXRXN_IN                   =>      GT0_GTXRXN_IN,
        GT0_GTXRXP_IN                   =>      GT0_GTXRXP_IN,
        GT0_RXCDRLOCK_OUT               =>      GT0_RXCDRLOCK_OUT,
        GT0_RXELECIDLE_OUT              =>      gt0_rxelecidle_i,
        -------- Receive Ports - RX Elastic Buffer and Phase Alignment Ports -------
        GT0_RXBUFRESET_IN               =>      GT0_RXBUFRESET_IN,
        GT0_RXBUFSTATUS_OUT             =>      GT0_RXBUFSTATUS_OUT,
        ------------------------ Receive Ports - RX PLL Ports ----------------------
        GT0_RXRESETDONE_OUT             =>      gt0_rxresetdone_i,
        ------------------------------- Transmit Ports -----------------------------
        GT0_TXUSERRDY_IN                =>      gt0_txuserrdy_i,
        ---------------- Transmit Ports - 8b10b Encoder Control Ports --------------
        GT0_TXCHARDISPMODE_IN           =>      GT0_TXCHARDISPMODE_IN,
        GT0_TXCHARDISPVAL_IN            =>      GT0_TXCHARDISPVAL_IN,
        GT0_TXCHARISK_IN                =>      GT0_TXCHARISK_IN,
        ------------ Transmit Ports - TX Buffer and Phase Alignment Ports ----------
        GT0_TXBUFSTATUS_OUT             =>      GT0_TXBUFSTATUS_OUT,
        ------------------ Transmit Ports - TX Data Path interface -----------------
        GT0_GTTXRESET_IN                =>      gt0_gttxreset_gt,
        GT0_TXDATA_IN                   =>      GT0_TXDATA_IN,
        GT0_TXOUTCLK_OUT                =>      GT0_TXOUTCLK_OUT,
        GT0_TXOUTCLKFABRIC_OUT          =>      GT0_TXOUTCLKFABRIC_OUT,
        GT0_TXOUTCLKPCS_OUT             =>      GT0_TXOUTCLKPCS_OUT,
        GT0_TXPCSRESET_IN               =>      gt0_txpcsreset_i,
        GT0_TXUSRCLK_IN                 =>      GT0_TXUSRCLK_IN,
        GT0_TXUSRCLK2_IN                =>      GT0_TXUSRCLK2_IN,
        ---------------- Transmit Ports - TX Driver and OOB signaling --------------
        GT0_GTXTXN_OUT                  =>      GT0_GTXTXN_OUT,
        GT0_GTXTXP_OUT                  =>      GT0_GTXTXP_OUT,
        ----------------------- Transmit Ports - TX PLL Ports ----------------------
        GT0_TXRESETDONE_OUT             =>      gt0_txresetdone_i



    );

    gt0_rxpcsreset_i                             <= tied_to_ground_i;
    gt0_txpcsreset_i                             <= tied_to_ground_i;





    GT0_CPLLLOCK_OUT                             <= gt0_cplllock_i;
    GT0_TXRESETDONE_OUT                          <= gt0_txresetdone_i;
    GT0_RXRESETDONE_OUT                          <= gt0_rxresetdone_i;
    GT0_RXELECIDLE_OUT                           <= gt0_rxelecidle_i;
    GT0_RXOUTCLK_OUT                             <= gt0_rxoutclk_i;

chipscope : if EXAMPLE_USE_CHIPSCOPE = 1 generate
    gt0_cpllreset_i                              <= GT0_CPLLRESET_IN;
    gt0_gttxreset_i                              <= GT0_GTTXRESET_IN;
    gt0_gtrxreset_i                              <= GT0_GTRXRESET_IN;
    gt0_txuserrdy_i                              <= GT0_TXUSERRDY_IN;
    gt0_rxuserrdy_i                              <= GT0_RXUSERRDY_IN;
end generate chipscope;

no_chipscope : if EXAMPLE_USE_CHIPSCOPE = 0 generate
       gt0_cpllreset_i <=   gt0_cpllreset_t ;
    gt0_cpllreset_i                              <= gt0_cpllreset_t;
    gt0_gttxreset_i                              <= gt0_gttxreset_t;
    gt0_gtrxreset_i                              <= gt0_gtrxreset_t;
    gt0_txuserrdy_i                              <= gt0_txuserrdy_t;
    gt0_rxuserrdy_i                              <= gt0_rxuserrdy_t;
end generate no_chipscope;


gt0_txresetfsm_i:  gig_eth_pcs_pma_v11_4_TX_STARTUP_FSM 

  generic map(
           GT_TYPE                  => "GTX", --GTX or GTH or GTP
           STABLE_CLOCK_PERIOD      => STABLE_CLOCK_PERIOD,           -- Period of the stable clock driving this state-machine, unit is [ns]
           RETRY_COUNTER_BITWIDTH   => 8, 
           TX_QPLL_USED             => FALSE ,                       -- the TX and RX Reset FSMs must
           RX_QPLL_USED             => FALSE,                        -- share these two generic values
           PHASE_ALIGNMENT_MANUAL   => FALSE                 -- Decision if a manual phase-alignment is necessary or the automatic 
                                                                     -- is enough. For single-lane applications the automatic alignment is 
                                                                     -- sufficient              
             )     
    port map ( 
        STABLE_CLOCK                    =>      SYSCLK_IN,
        TXUSERCLK                       =>      GT0_TXUSRCLK_IN,
        SOFT_RESET                      =>      SOFT_RESET_IN,
        QPLLREFCLKLOST                  =>      tied_to_ground_i,
        CPLLREFCLKLOST                  =>      gt0_cpllrefclklost_i,
        QPLLLOCK                        =>      tied_to_vcc_i,
        CPLLLOCK                        =>      gt0_cplllock_i,
        TXRESETDONE                     =>      gt0_txresetdone_sync,
        MMCM_LOCK                       =>      tied_to_vcc_i,
        GTTXRESET                       =>      gt0_gttxreset_t,
        MMCM_RESET                      =>      open,
        QPLL_RESET                      =>      open,
        CPLL_RESET                      =>      gt0_cpllreset_t,
        TX_FSM_RESET_DONE               =>      GT0_TX_FSM_RESET_DONE_OUT,
        TXUSERRDY                       =>      gt0_txuserrdy_t,
        RUN_PHALIGNMENT                 =>      open,
        RESET_PHALIGNMENT               =>      open,
        PHALIGNMENT_DONE                =>      tied_to_vcc_i,
        RETRY_COUNTER                   =>      open
           );






gt0_rxresetfsm_i:  gig_eth_pcs_pma_v11_4_RX_STARTUP_FSM 

  generic map(
           EXAMPLE_SIMULATION       => EXAMPLE_SIMULATION,
           GT_TYPE                  => "GTX", --GTX or GTH or GTP
           EQ_MODE                  => "DFE",
           STABLE_CLOCK_PERIOD      => STABLE_CLOCK_PERIOD,           --Period of the stable clock driving this state-machine, unit is [ns]
           RETRY_COUNTER_BITWIDTH   => 8, 
           TX_QPLL_USED             => FALSE ,                       -- the TX and RX Reset FSMs must
           RX_QPLL_USED             => FALSE,                        -- share these two generic values
           PHASE_ALIGNMENT_MANUAL   => FALSE                         -- Decision if a manual phase-alignment is necessary or the automatic 
                                                                     -- is enough. For single-lane applications the automatic alignment is 
                                                                     -- sufficient              
             )     
    port map ( 
        STABLE_CLOCK                    =>      SYSCLK_IN,
        RXUSERCLK                       =>      GT0_RXUSRCLK_IN,
        SOFT_RESET                      =>      SOFT_RESET_IN,
        QPLLREFCLKLOST                  =>      tied_to_ground_i,
        CPLLREFCLKLOST                  =>      gt0_cpllrefclklost_i,
        QPLLLOCK                        =>      tied_to_vcc_i,
        CPLLLOCK                        =>      gt0_cplllock_i,
        RXRESETDONE                     =>      gt0_rxresetdone_sync,
        MMCM_LOCK                       =>      tied_to_vcc_i,
        RECCLK_STABLE                   =>      gt0_recclk_stable_i,
        RECCLK_MONITOR_RESTART          =>      tied_to_ground_i,
        DATA_VALID                      =>      GT0_DATA_VALID_IN,
        TXUSERRDY                       =>      tied_to_vcc_i,
        GTRXRESET                       =>      gt0_gtrxreset_t,
        MMCM_RESET                      =>      open,
        QPLL_RESET                      =>      open,
        CPLL_RESET                      =>      open,
        RX_FSM_RESET_DONE               =>      GT0_RX_FSM_RESET_DONE_OUT,
        RXUSERRDY                       =>      gt0_rxuserrdy_t,
        RUN_PHALIGNMENT                 =>      open,
        RESET_PHALIGNMENT               =>      open,
        PHALIGNMENT_DONE                =>      tied_to_vcc_i,
        RXDFEAGCHOLD                    =>      gt0_rxdfeagchold_i,
        RXDFELFHOLD                     =>      gt0_rxdfelfhold_i,
        RXLPMLFHOLD                     =>      gt0_rxlpmlfhold_i,
        RXLPMHFHOLD                     =>      gt0_rxlpmhfhold_i,
        RETRY_COUNTER                   =>      open
           );




  cdrlock_timeout:process(SYSCLK_IN)
  begin
    if rising_edge(SYSCLK_IN) then
        if(gt0_gtrxreset_i = '1') then
          rx_cdrlocked       <= '0';
          rx_cdrlock_counter <=  0                        after DLY;
        elsif (rx_cdrlock_counter = WAIT_TIME_CDRLOCK) then
          rx_cdrlocked       <= '1';
          rx_cdrlock_counter <= rx_cdrlock_counter        after DLY;
        else
          rx_cdrlock_counter <= rx_cdrlock_counter + 1    after DLY;
        end if;
    end if;
  end process;

gt0_recclk_stable_i                          <= rx_cdrlocked;

end RTL;


