package prbs_package is   
	type tap_array 				is array (0 to 3) of integer;	
end prbs_package;

package body prbs_package is
end prbs_package;
